library IEEE;
use IEEE.STD_LOGIC_1644.all;

entity  is
	port (
	
	);
end ;

architecture  of  is

begin

end ;