--librerias

entity tb.MEMORY is
end tb.MEMORY;

architecture behavior of tb.MEMORY is
