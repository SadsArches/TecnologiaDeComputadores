-- Hola